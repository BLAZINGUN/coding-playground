module branch_unit (rs1_in,rs2_in,opcode_6_to_2_in,funct3_in,branch_taken_out);
    
    input [31:0] rs1_in,rs2_in;
    input [4:0] opcode_6_to_2_in;
    input [2:0] funct3_in;

    output branch_taken_out;
    

endmodule