package fifo_pkg;


    `include fifo_write_xtn.sv
    `include fifo_read_xtn.sv
    `include fifo_write_gen.sv
    `include fifo_read_gen.sv
    `include fifo_write_drv.sv
    `include fifo_read_drv.sv
    `include fifo_write_mon.sv
    `include fifo_read_mon.sv
    `include fifo_reference_model.sv
    `include fifo_sb.sv
    `include fifo_env.sv

endpackage