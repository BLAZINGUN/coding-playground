`timescale 10ns/10ps

module gray2bin
        (input [3:0] G, //gray code output
         output [3:0] bin   //binary input
        );


reg [3:0] bin;

always @ (G)

begin

assign bin[3] = G[3];
assign bin[2] = G[3] ^ G[2];
assign bin[1] = G[3] ^ G[2] ^ G[1];
assign bin[0] = G[3] ^ G[2] ^ G[1] ^ G[0];
end

endmodule
