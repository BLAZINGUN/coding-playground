module tb;
real pi;
integer a;
initial
begin
a=14;
$display(real'(a));
$display(pi);
end


endmodule
