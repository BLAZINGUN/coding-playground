module top;
	int n="a";
	int t;
	initial
		begin
			t=int'(13.5);//explicit casting 
		$display(t);
		$display(n);//implict casting

		end







endmodule
