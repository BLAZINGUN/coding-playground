module clock_generation();


endmodule