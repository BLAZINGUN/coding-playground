`timescale 10ns/10ps

module decoder_3x8_dataflow (
	input [2:0] a,
    output [7:0] d );

assign d[0] = (~a[2])&(~a[1])&(~a[0]);
assign d[1] = (~a[2])&(~a[1])&(a[0]);
assign d[2] = (~a[2])&(a[1])&(~a[0]);
assign d[3] = (~a[2])&(a[1])&(a[0]);
assign d[4] = (a[2])&(~a[1])&(~a[0]);
assign d[5] = (a[2])&(~a[1])&(a[0]);
assign d[6] = (a[2])&(a[1])&(~a[0]);
assign d[7] = (a[2])&(a[1])&(a[0]);

endmodule
