//when values need to be assigned between two different data type variables, ordinary assignment might not be valid and instead a system task called $cast should be used
//$cast can also be used as a function , but it returns 1 if the cast is legal

