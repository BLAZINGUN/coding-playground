module top();

class sub;

	int a;
endclass

/*class Base;
	int c;
	sub sbh= new;//sub class

endclass
Base bh1,bh2;
initial
	begin
		bh1=new;
		bh1.c=23;
		$display(bh1.c);
		bh1.sbh.a=34;
		$display(bh1.sbh.a);
		bh2 = new bh1;
		$display(bh1);
		$display(bh2);	
		$display(bh1.sbh);
		$display(bh2.sbh);	
			
	end

endmodule*/



/*module top();
int p,y;
	function  int num( int a);
		num=a+1;	
	endfunction

initial
	begin
	y=9;
	p=num(y);
	$display(p);
	end 
endmodule*/
