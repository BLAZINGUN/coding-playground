module top;

	int t ;
	initial
		begin
		t=int unsigned'(-13);
		$display(t);
		end





endmodule 
