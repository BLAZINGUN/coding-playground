module integer_file(clk_in,rst_in,rs_2_addr_in,rd_addr_in,wr_en_in,rd_in,rs_1_addr_in,rs_1_out,rs_2_out);

input clk_in,rst_in,wr_en_in;
input [31:0] rd_in;
input [4:0] rs_2_addr_in,rd_addr_in,rs_1_addr_in;

output [31:0] rs_1_out,rs_2_out;




















endmodule