module alu(op_1_in,op_2_in,opcode_in,result_out);

input [31:0] op_1_in,op_2_in;
input [3:0] opcode_in;

output [31:0] result_out;

endmodule