module ha(intr it);

assign 
